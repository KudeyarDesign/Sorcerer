-- Project Sorcerer - RISC-V core
--
-- Console Terminal for Avalon MM Bus and VGA output 
--

--
-- Copyright (C) 2017
-- Alexey Shistko     alexey@kudeyar.com
-- Andrei Safronov    andrei@kudeyar.com
--
-- This program is free software; you can redistribute it and/or
-- modify it under the terms of the GNU General Public License
-- as published by the Free Software Foundation; either version 2
-- of the License, or (at your option) any later version.
--
-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with this program; if not, write to the Free Software
-- Foundation, Inc., 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.STD_LOGIC_ARITH.all;			 
use IEEE.NUMERIC_STD.all;		 
use work.utils.all;

entity console_out is
	generic
	(
	  ROW_NUM: natural := 34;
		COL_NUM: natural := 80;
		BLINKED_CURSOR: natural range 0 to 1 := 0
	);
  port
  (
		reset: in std_logic;
		clk:   in std_logic;
		
		-- Avalon Slave
		avs_s1_chipselect: in std_logic;
		avs_s1_read: in std_logic;
		avs_s1_write: in std_logic;
		avs_s1_writedata: in std_logic_vector(7 downto 0);
		avs_s1_readdata: out std_logic_vector(7 downto 0);

--		sync: out std_logic;
		RED: out std_logic_vector(7 downto 0);
		GREEN: out std_logic_vector(7 downto 0);
		BLUE:  out std_logic_vector(7 downto 0);
		nRAMDAC_BLANK: out std_logic;
		nRAMDAC_SYNC: out std_logic;
		RAMDAC_CLK: out std_logic;
		HSYNC: out std_logic;
		VSYNC: out std_logic
	
--    DVI_D: out std_logic_vector(11 downto 0);
--	  DVI_DE: out std_logic;
--	  DVI_CLK: out std_logic	
  );	
end console_out;

architecture behaviour of console_out is	
  type color24 is record
    r: std_logic_vector(7 downto 0);
	 g: std_logic_vector(7 downto 0);
	 b: std_logic_vector(7 downto 0);
  end record;

  constant AMBER: color24 := (r => x"FF", g => x"7F", b => x"00");
  constant COLOR_FG: color24 := AMBER;
  
  constant FONT_WIDTH: natural := 8;
	constant FONT_HEIGHT: natural := 14; 
	constant FONT_W_BITS: natural := ceil_log2(FONT_WIDTH);
	constant FONT_H_BITS: natural := 4; -- port_bits(FONT_HEIGHT);
	
	constant FONT_SIZE: natural := 24576; 
  constant vga_font : std_logic_vector(0 to FONT_SIZE-1) :=
   "0001110111111000111111010101101100000000000000000000000000000000"  &   -- 0
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 64
   "0000000000000000000000000000000000000000000000010000000000000000"  &   -- 128
   "0000000000000000000000000000000000000000000000000000000001000000"  &   -- 192
   "1111111110001111111110111111111000000000000000000000000000000000"  &   -- 256
   "0000000000000000000000000000000000000000000000000000000000000001"  &   -- 320
   "0001101000010001010001100000100000000011010000110000100000000010"  &   -- 384
   "0000000000000000010101010101010110000000000010001010000001000000"  &   -- 448
   "1111111110001111111110111111111000000000000000000000000000000000"  &   -- 512
   "0000000000000000000000000000000000000000000000000000000000000001"  &   -- 576
   "1011111000110011011011100101100000000011011000110000100000100010"  &   -- 640
   "0000000000000000010101010101010110100100100010001010000000010000"  &   -- 704
   "1111111110001111111110111101111000000001000000000000000000000000"  &   -- 768
   "0000000000000000000000000000000010000000000000000000000000000000"  &   -- 832
   "1111011011101110011111000111000000000001011000110000000000100000"  &   -- 896
   "0101010101010101000000000000000001100100101000101000100000010000"  &   -- 960
   "1110000001011111000001111101100100000001000000000000000000000000"  &   -- 1024
   "0000000000000000000000000000000010000000000000000000000000000000"  &   -- 1088
   "0110111011111110000110100011110000000011011000110000100000100000"  &   -- 1152
   "0101010101010101010101010101010101000100010001101001000000100100"  &   -- 1216
   "1000000000000000000000000000000000000001000000000000000000000000"  &   -- 1280
   "0000000000000000000000000000000010000000000000000000000000000001"  &   -- 1344
   "0001101000010011010001100000110000000011011000110000100000000010"  &   -- 1408
   "0000000000000000010101010101010100000000010001000001000000100100"  &   -- 1472
   "1000000000000000000000000000000000000000000000000000000000000000"  &   -- 1536
   "0000000000000000000000000000000000000000000000000000000000000001"  &   -- 1600
   "0001001000000001010001000000000000000000010000110000000000000010"  &   -- 1664
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 1728
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 1792
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 1856
   "0000000000000000000000000000000000000000000000010000000000000000"  &   -- 1920
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 1984
   "1111111111111111111111111111111100000000000000000000010100000000"  &   -- 2048
   "0010111010011110101001111010000000100000100110000000000000000000"  &   -- 2112
   "0001001000000000110001000000001000000001010000100000000000000000"  &   -- 2176
   "0000000000000000000000000000000000000000000000000000000000001011"  &   -- 2240
   "1000000000000000000001000000000000000000000000001011011111000011"  &   -- 2304
   "1010111110111111111111111111010000100000100110000000000000000111"  &   -- 2368
   "0011111000110011110011101001101100000101101000000000001010101010"  &   -- 2432
   "0000000000000000010101010101010100111100000100010100011001011011"  &   -- 2496
   "0000000000000000000000000010000000100010010000001011011111000011"  &   -- 2560
   "1111111101101001111110000111010000100000100110000000100000000111"  &   -- 2624
   "0110110101110111100110101011101100011110101000001011101011101010"  &   -- 2688
   "0000000000000000010101010101010111111100001110111110111001010010"  &   -- 2752
   "0000000000000000000000000000000001101011010000001111011111000001"  &   -- 2816
   "1111111101101001111110000011011010001010010010000000100000001110"  &   -- 2880
   "1101001101000100111101001110011100011010000000001011101001000000"  &   -- 2944
   "0101010101010101000000000000000011110000111011101111110000110110"  &   -- 3008
   "0000001111010000111111000000001101000011100000001111111111001001"  &   -- 3072
   "1111111101100001111110000011011010001010011000000000000000011000"  &   -- 3136
   "1011111110111000111011101101110100011010101000001011101010101000"  &   -- 3200
   "0101010101010101010101010101010100101100111101110001101000111100"  &   -- 3264
   "0000000000000000000000000000000000100001100000001011111111001001"  &   -- 3328
   "1011011111010111111111111111010010001010001000000000000000010011"  &   -- 3392
   "0011110110111011010011101001100100001101101000000000001010101010"  &   -- 3456
   "0000000000000000010101010101010100011100000100110100011000001001"  &   -- 3520
   "1000000000000000000000000000000000100000000000000000010100000000"  &   -- 3584
   "0000011010010110000011111110000000000000000000000000000000010011"  &   -- 3648
   "0000000000000011000000001000000000000101000000000000001000001010"  &   -- 3712
   "0000000000000000000000000000000000010000000000000100010000000001"  &   -- 3776
   "1000000000000000000000000000000000000000000000000000000000000000"  &   -- 3840
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 3904
   "0000000000000000000000000000000000000000010000100000001000000000"  &   -- 3968
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 4032
   "1001111111101100111111011101111100000000000000001011011111000001"  &   -- 4096
   "1000000110010111010101111010000000000000000000000000000000000010"  &   -- 4160
   "0000001000000000000000001000000100000001010000100000001000001000"  &   -- 4224
   "1000000000000000000000000000000000110000000000000100010000011001"  &   -- 4288
   "0111111111011011000000110101101000001010000000001111011111000001"  &   -- 4352
   "1111111110011111111111111111000000100000100100000000000000000010"  &   -- 4416
   "0000001100000000100000001000001100011101001000001011001001101000"  &   -- 4480
   "1000000000000000010101010101010101111000001100111100111000011011"  &   -- 4544
   "0111111111001011000001110111101000101010000000000100000000000010"  &   -- 4608
   "0111111000001010101000000101001000100010100110000000100000000000"  &   -- 4672
   "0010010100000000100000000000001000011100101000101011000011100000"  &   -- 4736
   "1000000000000000010101010101010101001100011101111001101001100110"  &   -- 4800
   "1110001111010011000000100000111001101000110000000100100000001010"  &   -- 4864
   "0000000001100000000010000000001010000010010010000000100000011110"  &   -- 4928
   "0010011000000000000000000000000000100000110000100000001011001000"  &   -- 4992
   "1101010101010101000000000000000010010100010011001111010101100100"  &   -- 5056
   "1000001001000000111111000000010101001011110000000100100000001000"  &   -- 5120
   "0100100001110000000010000000011010001000011000000000000000011110"  &   -- 5184
   "0010011000000000100000000000000000010000111000101011001010101000"  &   -- 5248
   "1101010101010101010101010101010110111100101110011110111100011000"  &   -- 5312
   "0000000000000000000000000000000000101011000000001011101111000001"  &   -- 5376
   "1111111110010111111101111110011000001010001000000000000000000010"  &   -- 5440
   "0000000100000000100000001000000100010101001000001011000000100000"  &   -- 5504
   "1000000000000000010101010101010100111000101100110100111000011001"  &   -- 5568
   "0000000000000000000000000000000000100000000000001011001111000001"  &   -- 5632
   "1011011110000111111111111110000000000010000000000000000000000000"  &   -- 5696
   "0000000100000000000000001000000100001101000000000000001000001000"  &   -- 5760
   "1000000000000000000000000000000000000000000000100000000000000001"  &   -- 5824
   "1000000000000000000000000000000000000000000000000000000000000000"  &   -- 5888
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 5952
   "0000000000000000000000000000000000000000010000100000001000001000"  &   -- 6016
   "1000000000000000000000000000000000000000000000000000000000000000"  &   -- 6080
   "1001111111101100111111011101111100001000000000001010011011000001"  &   -- 6144
   "1101000110010111010101110010100000000000000000000000000000000000"  &   -- 6208
   "0000001111110000010000001111100100000000010000100000101000011000"  &   -- 6272
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 6336
   "0000000000010000000000000000000000011100001000001010011011000001"  &   -- 6400
   "1111111110011111111101111101101000100000100100000000000000000001"  &   -- 6464
   "0000001111110000111111101111111100111011000000000000101000011010"  &   -- 6528
   "0000000000000000010101010101010100000011000000000000000000000010"  &   -- 6592
   "0000000000000000000000000010001000010110101000000000100000001000"  &   -- 6656
   "0010111000001110101000001101001000100010100110000000100000000001"  &   -- 6720
   "1101100011111111101111100000011000111111011100101000100001100011"  &   -- 6784
   "0000000000000000010101010101010100000011000000000000000000000010"  &   -- 6848
   "1000000000010000000001000000000001101011100100000100100000001010"  &   -- 6912
   "0000000001110000000010000000000000000010000010000000100000011100"  &   -- 6976
   "1101101011111111001111100000001001100110001100001111101001111001"  &   -- 7040
   "0101010101010101000000000000000000000011000000000000000100000000"  &   -- 7104
   "1110001111000011111111100000010101010011011100000100100100110010"  &   -- 7168
   "0000000001110100000010001010010010001000000000000000000000011100"  &   -- 7232
   "1101101011111111001111101000001001100110001000001111101000111000"  &   -- 7296
   "0101010101010101010101010101010100000011000000001000000100000000"  &   -- 7360
   "0000000000000000000000000000000000111000011000011011100111110001"  &   -- 7424
   "1110100110000111111001111110011010001000000000000000000000000001"  &   -- 7488
   "0000000011111111111111101111111100100110011100100000100000000010"  &   -- 7552
   "0000000000000000010101010101010100000011000000001000000000000000"  &   -- 7616
   "0000000000000000000000000000000000001100000000011011000011000001"  &   -- 7680
   "1110100110000111111001110100001000000000000000000000000000000001"  &   -- 7744
   "0000000011110000110000001111110100000000001100000000101000001010"  &   -- 7808
   "0000000000000000000000000000000000000010000000000000000000000000"  &   -- 7872
   "1000000000000000000000000000000000000000000000000000000000000000"  &   -- 7936
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 8000
   "0000000000000000000000000000000000000000010000100000001000001000"  &   -- 8064
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 8128
   "1111111111101011111111110111101000010000000000001000011011000100"  &   -- 8192
   "1101000110010111010001110000000000000000000000101010111111100000"  &   -- 8256
   "0000001100000000011111101111100100101010010000100000111010001000"  &   -- 8320
   "0000000000000000000000001111111100000011000000000100000001111101"  &   -- 8384
   "1111110110100111111110111111010100011100000000001000111011001100"  &   -- 8448
   "1111111110011111111101110101100001111101110101111111111111100001"  &   -- 8512
   "1111111111110000111111111111111100111011100100000001111010011110"  &   -- 8576
   "0000000000000000010111111111111111111111111100001111111011111111"  &   -- 8640
   "1111110110110111111110111111010100011110101000000000100000001100"  &   -- 8704
   "0010111000011110101100001101100001111111110111010101100000100001"  &   -- 8768
   "1111110011110000110000010000011000011001110100100011000011010111"  &   -- 8832
   "0000000000000000011111111111111111111100111111111011111010000010"  &   -- 8896
   "1111110110100111111110111111011101011010101100000100000100000100"  &   -- 8960
   "1000000001110110000010001010000001111111011010111111100000111100"  &   -- 9024
   "0010011000001111000000001000000001101101100000000110001011001001"  &   -- 9088
   "0101010101010101001010101010101011111110111111111111111010000010"  &   -- 9152
   "0000001001100100000001011111000001010010011100010110100100110111"  &   -- 9216
   "1000000001100100000010001010010001111100111001111011110000111100"  &   -- 9280
   "1111111000001111000000011000000001001101100100000101011010011100"  &   -- 9344
   "0101010101010101011111111111111111111110111111111111111011111010"  &   -- 9408
   "0000000000000000000000000000000000010100010000011011100011110111"  &   -- 9472
   "1110100010000111111001110100010000111101101101111111111111100001"  &   -- 9536
   "1111110011110000111111111111111100100011100100100001110010011110"  &   -- 9600
   "0000000000000000011111111111111100000001111100001111111011111101"  &   -- 9664
   "1000000000000000000000000000000000010100000000001001000011000100"  &   -- 9728
   "1110100010000111111001110100000000000001000100000100001111100001"  &   -- 9792
   "0000000011110000111111101111111100100010000000000000101010001010"  &   -- 9856
   "0000000000000000001100110011001100000011000000001000000010000101"  &   -- 9920
   "1000000000000000000000000000000000000000000000000000000000000000"  &   -- 9984
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 10048
   "0000000000000000000000000000000000000000010000100000001000001000"  &   -- 10112
   "0000000000000000001100110011001100000010000000000000000000000000"  &   -- 10176
   "1000000000000000000000000000000000000000001001001000111000001000"  &   -- 10240
   "1101000110010111010001110000000000011111000001010101011101100000"  &   -- 10304
   "1111111100000000111111101111100100110011110100100000010010001100"  &   -- 10368
   "0000000011111111000000000000000000000001111100001011111011111101"  &   -- 10432
   "1000000000000000000000000000000000010010001101001000111011001000"  &   -- 10496
   "1111111110011111111001110001000000111111100101111111011111010001"  &   -- 10560
   "1111111111110000111111101111111100111111101111000110011001101100"  &   -- 10624
   "0000000011111111010111110000000000000001111100001111111111111111"  &   -- 10688
   "1000000000000000000000000000000000011010101101000001011111000000"  &   -- 10752
   "0010111010011000101100001111100000100010100111101010100010010001"  &   -- 10816
   "0000001011110000110000010000011000011100011011100111001001110010"  &   -- 10880
   "0000000011111111011111110000000000000000000000000100000100000010"  &   -- 10944
   "0000000000000000000000000000000001001010101101011111011111000001"  &   -- 11008
   "1010011011110110101110011110100000000010110011000000100000011000"  &   -- 11072
   "0000001000001111110000011000000000110100001111100111001101111110"  &   -- 11136
   "0111111111111111001000000000000000000010000011110000000100000000"  &   -- 11200
   "0000000000000000000000000000000001011100011101010111111011000001"  &   -- 11264
   "1010011011100000101110001100010001001011011101000100010010101100"  &   -- 11328
   "0000001000001111000000010000000100000100001111100111111111101110"  &   -- 11392
   "0111111111111111010011001100110011111110000011110000000111111010"  &   -- 11456
   "1000000000000000000000000000000000010100011101001001111011000010"  &   -- 11520
   "1110111010000111111001110100010001111111101101111111011111100101"  &   -- 11584
   "1111111000000000111111101111111100000101101011000110110010110010"  &   -- 11648
   "0011001100110011010011001100110011111100111100001111111111111111"  &   -- 11712
   "1000000000000000000000000000000000000010001101001000000001000010"  &   -- 11776
   "1100100010000111010001110000000000110101100001111011001101000101"  &   -- 11840
   "1111111000000000111111101111111000000101101011000100001000010100"  &   -- 11904
   "0011001100110011000000000000000000000010111100001111111110000101"  &   -- 11968
   "1000000000000000000000000000000000000000000000000000000000000000"  &   -- 12032
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 12096
   "0000000000000000000000000000000000000000010000100000001000000000"  &   -- 12160
   "0011001100110011000000000000000000000010000000000000000000000000"  &   -- 12224
   "1000000000000000000000000000000000000010000000001000101010000100"  &   -- 12288
   "1101000110010111010001110000000000011101000001010100011101000000"  &   -- 12352
   "1111111100000000011111101111100100101001010000100000010000001100"  &   -- 12416
   "0000000000000000000000001111111100000001111100001011111011111101"  &   -- 12480
   "1000000000000000000000000000000000010010000000001000101010001100"  &   -- 12544
   "1111111110011111111001110011000001111101100101111111011101000000"  &   -- 12608
   "1111111111110000111111101111101100111011100100000000010000011100"  &   -- 12672
   "0000000000000000010111111111111111111111111100001111111011111111"  &   -- 12736
   "1000000000000000000000000000000000010010101000010010100100001100"  &   -- 12800
   "0110111000001000101000011011000001100110100110101011100010000001"  &   -- 12864
   "0000000011110000100000011000011000011010110100100000100000010001"  &   -- 12928
   "0000000000000000011111111111111111111110111100000100000000000010"  &   -- 12992
   "0111100001111100000100111100000001001110101100010110100100000101"  &   -- 13056
   "1100000001110010001010011100100001000110010111000001100110111101"  &   -- 13120
   "0000001011111111010000011000010001101110100000000100101110001111"  &   -- 13184
   "0000111100001111011100001111000011111110111111110000000010000000"  &   -- 13248
   "0000111111111111111101010010111101011110011100000100100000000111"  &   -- 13312
   "1100000101110010001110011100110001001100011100000100010010111101"  &   -- 13376
   "0000001011111111010000010000010001001110000100000100111110011110"  &   -- 13440
   "0000111100001111011111111111111111111110111111110000000011111010"  &   -- 13504
   "1000110011111111011110010011111100011010010000001001111011000110"  &   -- 13568
   "1110100110000111010101110000010001101101101001111100011101000001"  &   -- 13632
   "1111110111110000111111101111111100000011010110100000010000010100"  &   -- 13696
   "0000000000000000011111111111111111111110111100001111111011111111"  &   -- 13760
   "1000110011111111000010010011111100000010000000001001111011000100"  &   -- 13824
   "1110100110000111010001110000000000100101100001111000001101000000"  &   -- 13888
   "1111110100000000111111101111101100000001000010000000001000000100"  &   -- 13952
   "0000000000000000001100110011001100000010111100001111111010000101"  &   -- 14016
   "1111101011111000000001101101111100000000000000000000000000000000"  &   -- 14080
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 14144
   "0000000000000000000000000000000000000000010000100000001000000000"  &   -- 14208
   "0000000000000000001100110011001100000010000000000000000000000000"  &   -- 14272
   "1000000000000000000000000000000000001010000000001000001010000000"  &   -- 14336
   "1101000110110111010001010010000001011101000001010100010101000000"  &   -- 14400
   "1111111000000000011111101111100100100000010000100000010000011100"  &   -- 14464
   "0000000000000000100000000000000011111111111100001011111011111101"  &   -- 14528
   "1000000000000000000000000000000000011010001000011010001010000000"  &   -- 14592
   "1111111110011111111001111011000001111101100101111110011101000000"  &   -- 14656
   "1111111111110000111111111111101100111001000000000000110000011100"  &   -- 14720
   "0000000000000000100011110000111111111111111100001111111011111111"  &   -- 14784
   "1000000000000000000000000000000000010100101000010010000100001000"  &   -- 14848
   "0010111000001000101000111001000000100010100110101010101010100000"  &   -- 14912
   "1111110111110000100000011000001000011101000100100000100010000001"  &   -- 14976
   "0000000000000000100011110000111100000000000000000100000010000010"  &   -- 15040
   "1100010010101110011000011110111101001100100100000100000100001010"  &   -- 15104
   "1000000001100000000010000100000000000010010011000001100110111101"  &   -- 15168
   "1111111000001111000000000000011001100101110100000100001010011111"  &   -- 15232
   "0000111100001111100000000000000000000010000011110000000110000000"  &   -- 15296
   "1011001100000000100011101101000001010010011110000100100000110010"  &   -- 15360
   "1000000001110010001010111100110001001000011100000101011011011101"  &   -- 15424
   "1111111000001111010000010000011001000101110000000100011000011110"  &   -- 15488
   "0000111100001111100011110000111111111110000011110000000101111111"  &   -- 15552
   "1000100001010001010000000000000000011010011010001001111011110000"  &   -- 15616
   "1110100110010111011101111000110001101001101101111101011101000000"  &   -- 15680
   "1111110100000000111111111111101100110111100110100000010000000000"  &   -- 15744
   "0000000000000000100011110000111111111101000000001111111011111111"  &   -- 15808
   "1011001000000000001111100100000000001000000000001001011011000000"  &   -- 15872
   "0110100110001111010101010010000000100001100001111000000101000000"  &   -- 15936
   "1111110100000000111111101111100100110010000110000000101000000000"  &   -- 16000
   "0000000000000000100000000000000000000001000000001111111010000101"  &   -- 16064
   "1100010000000110000000011110000000000000000000000000000000000000"  &   -- 16128
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 16192
   "0000000000000000000000000000000000000000010000100000001000001000"  &   -- 16256
   "0000000000000000100000000000000000000000000000000000000000000000"  &   -- 16320
   "1000000000000000000000000000000000010010000000011011011011000000"  &   -- 16384
   "1100000110110111010101011010000001011100000001010001010100000000"  &   -- 16448
   "1111111000000000011111101111100100010010110000100000110000001100"  &   -- 16512
   "0000000000000000000000000000000011111110111100001011111011111000"  &   -- 16576
   "1000000000000000000000000000000000011110000000011011011011000000"  &   -- 16640
   "1111111110111111111101011011000001111101100101111111010111100000"  &   -- 16704
   "1111111011110000111111101111101100111010100000000000110010001101"  &   -- 16768
   "0000000000000000000011110000111111111111111100001111111011111111"  &   -- 16832
   "1000000000000000000000000000000000011100000000000000000100000010"  &   -- 16896
   "0011111000001000101000100001000000100011100110101110101111100000"  &   -- 16960
   "0000000111110000100000000000001001111000000000000000000010000001"  &   -- 17024
   "0000000000000000000011110000111100000001000000000100000010000111"  &   -- 17088
   "0100010000101110000010011110000000011000110000100100000100001011"  &   -- 17152
   "0000000001100000010010100100000001000011010010001100101101011101"  &   -- 17216
   "0000001100001111000000000000010101110100000000000000001000001110"  &   -- 17280
   "0000111100001111000000000000000011111111000011110000000100000111"  &   -- 17344
   "0100001110101100100011010011111100011010110010100100100000111001"  &   -- 17408
   "0000100001100010000010100100010001001001011000001100011110011101"  &   -- 17472
   "0000001100001111100000000000010001100101000000000000011000001110"  &   -- 17536
   "0000111100001111000011110000111111111111000011110000000101111010"  &   -- 17600
   "1111101011111101011111111110111100011110000010001011111011110000"  &   -- 17664
   "0111110110011111011101011010110001111101101101111101010111000000"  &   -- 17728
   "1111110111110000111111101111100101110011100010000000110000001000"  &   -- 17792
   "0000000000000000000011110000111111111101111100001111111011111101"  &   -- 17856
   "1100000010000100000010010010111100010100000000001011011011000000"  &   -- 17920
   "0111010110011111011101011010100000110101100101110001000101100000"  &   -- 17984
   "1111110011110000011111101111100100011010100010000000101010001100"  &   -- 18048
   "0000000000000000000000000000000000000010111100001111111010000101"  &   -- 18112
   "1100010000000110000000001110000000000000000000000000000000000000"  &   -- 18176
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 18240
   "0000000000000000000000000000000000000000010000100000001000001000"  &   -- 18304
   "0000000000000000000000000000000000000010000000000000000000000000"  &   -- 18368
   "1000000000000000000000000000000000000100000000000010000000000000"  &   -- 18432
   "0110111010011110101000011010000000100000101111000010000010100000"  &   -- 18496
   "1111111011110000110000001000001110000001000000000000110010000001"  &   -- 18560
   "0000000000000000000000000000000000000000000000000000000010000000"  &   -- 18624
   "1000000000000000000000000000000000010110000000001111011011000010"  &   -- 18688
   "1110111110111111111101011011010001111110111111111011010110100100"  &   -- 18752
   "1111111011110000111111101111101100010011110000100100110010001101"  &   -- 18816
   "0000000000000000000011110000111111111110111100001111111011111010"  &   -- 18880
   "1000000000000000000000000000000000010010010000001111011111000010"  &   -- 18944
   "1011111101101001111111000111010001111110110110111011010100100101"  &   -- 19008
   "0000000011111111101111101111111001011010110000100100110010001110"  &   -- 19072
   "0000000000000000000011110000111111111110111111111111111011111010"  &   -- 19136
   "0100010000101110000000011110000001001010010000101111011111000001"  &   -- 19200
   "1011111101101001110111100111010001111110010010010011111000101101"  &   -- 19264
   "0000001111111111101111101111111101101110110000100100111010000010"  &   -- 19328
   "0000111100001111000000000000000011111111111111111011111011111000"  &   -- 19392
   "0011001100000000101001000001000001010000100010101111111011011001"  &   -- 19456
   "1011110101001001010111000111010000111110011010010101100100111001"  &   -- 19520
   "0000001111111111101111101111110101011110110000100100101010001110"  &   -- 19584
   "0000111100001111000011110000111100000011111111111011111010000000"  &   -- 19648
   "1000100001010001010000100000000000010110100010001111111011011000"  &   -- 19712
   "1111010111011111011111011111010001111101111111110101110111110001"  &   -- 19776
   "1111111011111111011111101111110101011011110000100100110010001111"  &   -- 19840
   "0000000000000000000011110000111111111110111111111111111011111101"  &   -- 19904
   "1011011000000100000111001000000000000110000000000110000000000000"  &   -- 19968
   "1100010010011110001000011010000001001001110101100000010011110000"  &   -- 20032
   "1111111011110000010000000000000010000001010000100100111010001001"  &   -- 20096
   "0000000000000000000000000000000011111110000000000100000001111101"  &   -- 20160
   "1100010010000010000000011110111100000000000000000000000000000000"  &   -- 20224
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 20288
   "0000000000000000000000000000000000000000000000000000001000000000"  &   -- 20352
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 20416
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 20480
   "0000000000000000000000000000000000000001001000000000000001000000"  &   -- 20544
   "0000000100000000000000000000000110000001000000000000010000000001"  &   -- 20608
   "0000000000000000000000000000000000000000000000000000000000000101"  &   -- 20672
   "1000000000000000000000000000000000000000000000000000000000000000"  &   -- 20736
   "0000000000000000000000000000000000000001001000001000000001000000"  &   -- 20800
   "0000000100000000000000000000000010000001000000000000010000000001"  &   -- 20864
   "0000000000000000000011110000111100000001000000000000000000000111"  &   -- 20928
   "1000000000000000000000000000000000000000000000000000000000000000"  &   -- 20992
   "0000000000000000000000000000000000000000000000001000000000000000"  &   -- 21056
   "0000000000000000000000000000000011000000000000000000000000000000"  &   -- 21120
   "0000000000000000000011110000111100000001000000000000000000000010"  &   -- 21184
   "1111000010101100011100011110111101000000000010000000000000010000"  &   -- 21248
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 21312
   "0000000000000000000000000000000011000000000000000000000000000000"  &   -- 21376
   "0000111100001111000000000000000000000000000000000000000000000000"  &   -- 21440
   "1000011110000011111101010000111101000000000010000000000000010000"  &   -- 21504
   "0000000000000000000000000000000000000000001000000100000000000000"  &   -- 21568
   "0000000100000000000000000000000011000000000000000000000000000000"  &   -- 21632
   "0000111100001111000011110000111100000001000000000000000000000000"  &   -- 21696
   "1000110111010011111100110001111100000000000000000000000000000000"  &   -- 21760
   "0000000000000000010000000000000000000001001000000100000001000000"  &   -- 21824
   "0000000100000000000000000000000011000001000000000000000000000001"  &   -- 21888
   "0000000000000000000011110000111100000001000000000000000000000101"  &   -- 21952
   "1000010110000011111010010001111100000000000000000000000000000000"  &   -- 22016
   "0000000000000000010000000000000000000001000000000000000001000000"  &   -- 22080
   "0000000000000000000000000000000010000001000000000000000000000001"  &   -- 22144
   "0000000000000000000000000000000000000000000000000000000000000101"  &   -- 22208
   "0111001100000100110001001111000000000000000000000000000000000000"  &   -- 22272
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 22336
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 22400
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 22464
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 22528
   "0000000000000000000000000000000100000000000000001000000000000000"  &   -- 22592
   "0000000000000000000000000000000000000000000000000000010000000000"  &   -- 22656
   "0000000000000000000000000000000000000000000000000000000000000010"  &   -- 22720
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 22784
   "0000000000000000000000000000000100000001001000001000000001000000"  &   -- 22848
   "0000000000000000000000000000000000000001000000000000010000000001"  &   -- 22912
   "0000000000000000000011110000111100000000000000000000000000000111"  &   -- 22976
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 23040
   "0000000000000000000000000000000100000001001000001000000001000000"  &   -- 23104
   "0000000100000000000000000000000000000001000000000000000000000001"  &   -- 23168
   "0000000000000000000011110000111100000001000000000000000000000111"  &   -- 23232
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 23296
   "0000000000000000000000000000000100000001001000001100000001000000"  &   -- 23360
   "0000000100000000000000000000000001000001000000000000000000000001"  &   -- 23424
   "0000111100001111000000000000000000000001000000000000000000000111"  &   -- 23488
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 23552
   "0000000000000000000000000000000100000001001000000100000001000000"  &   -- 23616
   "0000000100000000000000000000000001000001000000000000000000000001"  &   -- 23680
   "0000111100001111000011110000111100000001000000000000000000000101"  &   -- 23744
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 23808
   "0000000000000000000000000000000100000001000000000100000001000000"  &   -- 23872
   "0000000000000000000000000000000000000001000000000000000000000001"  &   -- 23936
   "0000000000000000000011110000111100000000000000000000000000000101"  &   -- 24000
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 24064
   "0000000000000000000000000000000100000000000000000100000000000000"  &   -- 24128
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 24192
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 24256
   "0000010000000000000000000000000000000000000000000000000000000000"  &   -- 24320
   "0000000000000000000000000000000100000000000000000000000000000000"  &   -- 24384
   "0000000000000000000000000000000000000000000000000000000000000000"  &   -- 24448
   "0000000000000000000000000000000000000000000000000000000000000000"   -- 24512
;

  type font_rom_type is array (0 to FONT_SIZE/8-1) of std_logic_vector(7 downto 0);
	function initFont(f: std_logic_vector(0 to FONT_SIZE-1)) return font_rom_type is
	  variable v: font_rom_type;
		variable d: std_logic_vector(7 downto 0);
	begin
		for i in 0 to FONT_SIZE/8-1 loop
			d := (others => '0');
			for j in 0 to 7 loop
				d(j) := f(i*8 + j);
			end loop;
			v(i) := d;
		end loop;	
		return v;
	end function initFont;	
	
	signal font_rom: font_rom_type := initFont(vga_font); 

--  signal RED: std_logic_vector(7 downto 0);
--  signal GREEN: std_logic_vector(7 downto 0);
--  signal BLUE:  std_logic_vector(7 downto 0);
--  signal nRAMDAC_BLANK: std_logic;
--  signal nRAMDAC_SYNC: std_logic;
--  signal RAMDAC_CLK: std_logic;

	type VGA_timings is 
	record
		h_polarity: boolean;
	  h_visible_area: natural;
		h_front_porch: natural;
		h_sync_pulse: natural;
		h_back_porch: natural;
		whole_line: natural;	
		v_polarity: boolean;
	  v_visible_area: natural;
		v_front_porch: natural;
		v_sync_pulse: natural;
		v_back_porch: natural;
		whole_frame: natural;
	end record;
	
	-- 640 x 350 x 70 Hz , f = 25.175 Mhz
	constant VGA_640x350x70: VGA_timings :=
	(			
	  h_polarity => true,     -- positive
	  h_visible_area => 640,	-- 25.422045680238 us
		h_front_porch => 16,		-- 0.63555114200596 us
		h_sync_pulse => 96,			-- 3.8133068520357 us 
		h_back_porch => 48,	  	-- 1.9066534260179 us
		whole_line => 800,	 		-- 31.777557100298 us
		v_polarity => false,    -- negative
		v_visible_area => 350,	-- 11.122144985104 ms
		v_front_porch => 37,		-- 1.175769612711 ms
		v_sync_pulse => 2,			-- 0.063555114200596 ms
		v_back_porch => 60,			-- 1.9066534260179 ms
		whole_frame => 449			-- 14.268123138034 ms
	);
	
	-- 512 x 256 x 70 Hz , f = 25.175 Mhz
	constant BK_512x256x70: VGA_timings :=
	(			
	  h_polarity => true,     -- positive
	  h_visible_area => 512,	-- 
		h_front_porch => 80,		-- 
		h_sync_pulse => 96,			-- 
		h_back_porch => 112,	  -- 
		whole_line => 800,	 		-- 
		v_polarity => false,    -- negative
		v_visible_area => 256,	-- 
		v_front_porch => 84,		-- 
		v_sync_pulse => 2,			-- 
		v_back_porch => 107,			-- 
		whole_frame => 449			-- 
	);	
	
	-- 640 x 350 x 85 Hz , f = 31.5 Mhz
	constant VESA_640x350x85: VGA_timings :=
	(			
	  h_polarity => true,     -- positive
	  h_visible_area => 640,	-- 20.31746031746 us
		h_front_porch => 32,		-- 1.015873015873 us
		h_sync_pulse => 64,			-- 2.031746031746 us 
		h_back_porch => 96,	  	-- 3.047619047619 us
		whole_line => 832,	 		-- 26.412698412698 us
		v_polarity => false,    -- negative
		v_visible_area => 350,	-- 9.2444444444444 ms
		v_front_porch => 32,		-- 0.84520634920635 ms
		v_sync_pulse => 3,			-- 0.079238095238095 ms
		v_back_porch => 60,			-- 1.5847619047619 ms
		whole_frame => 445			-- 11.753650793651 ms
	);	
	
		-- 640 x 480 x 60 Hz , f = 25.175 Mhz	Industry standard timing
	constant VGA_640x480x60: VGA_timings :=
	(			
	  h_polarity => false,    -- negative
	  h_visible_area => 640,	-- 25.422045680238 us
		h_front_porch => 16,		-- 0.63555114200596 us
		h_sync_pulse => 96,			-- 3.8133068520357 us 
		h_back_porch => 48,		  -- 1.9066534260179 us
		whole_line => 800,	 		-- 31.777557100298 us
		v_polarity => false,    -- negative
		v_visible_area => 480,	-- 15.253227408143 ms
		v_front_porch => 10,		-- 0.31777557100298 ms
		v_sync_pulse => 2,			-- 0.063555114200596 ms
		v_back_porch => 33,			-- 1.0486593843098 ms
		whole_frame => 525			-- 16.683217477656 ms
	);
	
	-- 640 x 480 x 73 Hz , f = 31.5 Mhz
	constant VGA_640x480x73: VGA_timings :=
	(			
	  h_polarity => false,    -- negative
	  h_visible_area => 640,	-- 20.31746031746 us
		h_front_porch => 24,		-- 0.76190476190476 us
		h_sync_pulse => 40,			-- 1.2698412698413 us 
		h_back_porch => 128,		-- 4.0634920634921 us
		whole_line => 832,	 		-- 26.412698412698 us
		v_polarity => false,    -- negative
		v_visible_area => 480,	-- 12.678095238095 ms
		v_front_porch => 9,			-- 0.23771428571429 ms
		v_sync_pulse => 2,			-- 0.052825396825397 ms
		v_back_porch => 29,			-- 0.76596825396825 ms
		whole_frame => 520			-- 13.734603174603 ms
	);		
	
	-- 640 x 480 x 75 Hz , f = 31.5 Mhz
	constant VESA_640x480x75: VGA_timings :=
	(			
	  h_polarity => false,    -- negative
	  h_visible_area => 640,	-- 20.31746031746 us
		h_front_porch => 16,		-- 0.50793650793651 us
		h_sync_pulse => 64,			-- 2.031746031746 us 
		h_back_porch => 120,		-- 3.8095238095238 us
		whole_line => 840,	 		-- 26.666666666667 us
		v_polarity => false,    -- negative
		v_visible_area => 480,	-- 12.8 ms
		v_front_porch => 1,			-- 0.026666666666667 ms
		v_sync_pulse => 3,			-- 0.08 ms
		v_back_porch => 16,			-- 0.42666666666667 ms
		whole_frame => 500			-- 13.333333333333 ms
	);	
	
	-- 768 x 576 x 75 Hz , f = 45.51 Mhz
	constant VESA_768x576x75: VGA_timings :=
	(			
	  h_polarity => false,    -- negative
	  h_visible_area => 768,	-- 16.875411997363 us
		h_front_porch => 40,		-- 0.878927708196 us
		h_sync_pulse => 80,			-- 1.757855416392 us 
		h_back_porch => 120,		-- 2.636783124588 us
		whole_line => 1008,	 		-- 22.148978246539 us
		v_polarity => true,     -- positive
		v_visible_area => 576,	-- 12.757811470007 ms
		v_front_porch => 1,			-- 0.022148978246539 ms
		v_sync_pulse => 3,			-- 0.066446934739618 ms
		v_back_porch => 22,			-- 0.48727752142386 ms
		whole_frame => 602			-- 13.333684904417 ms
	);	
	
	-- 800 x 600 x 72 Hz , f = 50.0 Mhz
	constant VGA_640x480x72: VGA_timings :=
	(										 
	  h_polarity => true,		  -- pisitive
	  h_visible_area => 800,	-- 16 us
		h_front_porch => 56,		-- 1.12 us
		h_sync_pulse => 120,		-- 2.4 us
		h_back_porch => 64,			-- 1.28 us
		whole_line => 1040,			-- 20.8 us
		v_polarity => true,		  -- positive
		v_visible_area => 600,	-- 12.48 ms
		v_front_porch => 37,		-- 0.7696 ms
		v_sync_pulse => 6,			-- 0.1248 ms
		v_back_porch => 23,			-- 0.4784 ms
		whole_frame => 666      -- 13.8528 ms
	);	
	
  type internal_timings is 
  record
		h_sync_inv: std_logic;
  	h_sync_end: std_logic_vector(10 downto 0);
	  h_blank_start: std_logic_vector(10 downto 0);
	  h_blank_end: std_logic_vector(10 downto 0);
	  h_size: std_logic_vector(10 downto 0);
		v_sync_inv: std_logic;
    v_sync_end: std_logic_vector(10 downto 0);
	  v_blank_start: std_logic_vector(10 downto 0);
	  v_blank_end: std_logic_vector(10 downto 0);
	  v_size: std_logic_vector(10 downto 0);	
	end record;

	function convert_timings(t: VGA_timings) return internal_timings is
	  variable v: internal_timings;
		variable v_delta: natural;
	begin																	
		assert t.h_visible_area + t.h_front_porch+ t.h_sync_pulse+ t.h_back_porch = t.whole_line 
		  report "Invalid horizontal timings" severity error;	
		assert t.v_visible_area + t.v_front_porch+ t.v_sync_pulse+ t.v_back_porch = t.whole_frame 
		  report "Invalid vertical timings" severity error;		
		if t.h_polarity then
			v.h_sync_inv := '0';
		else
			v.h_sync_inv := '1';
		end if;	
		v.h_sync_end := conv_std_logic_vector(t.h_sync_pulse- 1, 11);
		v.h_blank_start := conv_std_logic_vector(t.whole_line- t.h_front_porch- 1, 11);
		v.h_blank_end := conv_std_logic_vector(t.h_sync_pulse+ t.h_back_porch- 1, 11);
	  v.h_size := conv_std_logic_vector(t.whole_line- 1, 11);
		if t.v_polarity then
			v.v_sync_inv := '0';
		else
			v.v_sync_inv := '1';
		end if;		
		v.v_sync_end := conv_std_logic_vector(t.v_sync_pulse- 1, 11);
		v_delta := t.v_visible_area - ROW_NUM * FONT_HEIGHT;
		v.v_blank_start := conv_std_logic_vector(t.whole_frame- t.v_front_porch- 1 - v_delta, 11);
		v.v_blank_end := conv_std_logic_vector(t.v_sync_pulse+ t.v_back_porch- 1, 11);
		v.v_size := conv_std_logic_vector(t.whole_frame- 1, 11);
		return v;
	end function;	

	signal clk_en: std_logic;
	
	signal tms: internal_timings;

	signal blank: std_logic;
	signal blank_del, blank_del2, blank_del3: std_logic;
	
	constant X_BITS: natural := 7;
	constant Y_BITS: natural := 6;
	constant CHAR_RAM_SIZE: natural := ROW_NUM* COL_NUM;
	constant CHAR_RAM_BITS: natural := Y_BITS + X_BITS;

	type char_ram_type is array (0 to CHAR_RAM_SIZE) of std_logic_vector(7 downto 0);
	signal char_ram: char_ram_type;
	signal char_ram_q: std_logic_vector(7 downto 0);
	
	type char_ram_cmd_type is record
		rd_address: std_logic_vector(CHAR_RAM_BITS-1 downto 0);		
		wr_address: std_logic_vector(CHAR_RAM_BITS-1 downto 0);
		wr_data: std_logic_vector(7 downto 0);
		wr: std_logic;
	end record;	
	signal char_ram_cmd: char_ram_cmd_type;

	signal font_rom_address: std_logic_vector(11 downto 0);
	signal font_rom_q: std_logic_vector(7 downto 0);
	
	type state_type is (st_clear_screen, st_clear_row, st_idle, st_tab);
	type display_regs_type is record	
		state: state_type;
		
		display_clk_cnt: std_logic_vector(0 downto 0);
	  hcnt: std_logic_vector(10 downto 0);
	  vcnt: std_logic_vector(10 downto 0);
	  hblank: std_logic;
	  hsync: std_logic;
	  vblank: std_logic;
	  vsync: std_logic;			
		
		cursor_x: std_logic_vector(X_BITS- 1 downto 0);
		cursor_y: std_logic_vector(Y_BITS-1 downto 0);
		rd_ptr_x: std_logic_vector(X_BITS-1 downto 0);
		rd_ptr_y: std_logic_vector(Y_BITS-1 downto 0);
		scroll_y: std_logic_vector(Y_BITS-1 downto 0);
		font_row: std_logic_vector(FONT_H_BITS-1 downto 0);
		font_col: std_logic_vector(FONT_W_BITS-1 downto 0);
		font_lsb: std_logic_vector(2 downto 0);
		
	  rcolor: std_logic_vector(7 downto 0);
	  gcolor: std_logic_vector(7 downto 0);
	  bcolor: std_logic_vector(7 downto 0);			
		
    cursor_cnt: std_logic_vector(5 downto 0);	
		
    sym: std_logic_vector(7 downto 0);
	  sym_rdy: std_logic;		
	end record; 
	
	signal r, next_r: display_regs_type;
	
	function get_address(x: std_logic_vector(X_BITS- 1 downto 0); 
	    y: std_logic_vector(Y_BITS-1 downto 0); scroll_y: std_logic_vector(Y_BITS-1 downto 0)) 
	    return std_logic_vector is
		variable y1, y2: std_logic_vector(Y_BITS downto 0);	
		variable ya: std_logic_vector(Y_BITS-1 downto 0);
		variable address, da: std_logic_vector(CHAR_RAM_BITS-1 downto 0);
	begin	 	
		da := (others => '0');
		address := (others => '0');
		y1 := ('0' & y) + ('0' & scroll_y);
		y2 := y1 - CONV_STD_LOGIC_VECTOR(ROW_NUM, Y_BITS+ 1);
		if y2(Y_BITS) = '1' then
			ya := y1(Y_BITS-1 downto 0);
		else	
			ya := y2(Y_BITS-1 downto 0);
		end if;	
		case COL_NUM is	
			when 64 =>
			  address(Y_BITS+5 downto 6) := ya;
			when 80 =>
			  address(Y_BITS+5 downto 6) := ya;
				da(Y_BITS+3 downto 4) := ya;
				address := address + da;
			when others => null;  -- TODO
		end case;	
		address := address + x;
	  return address;	
	end function get_address;	
begin	
	tms <= convert_timings(VGA_640x480x60);
--	tms <= convert_timings(VGA_640x350x70);
	
	
	next_state_proc: process(r,	clk_en,
    	avs_s1_chipselect, avs_s1_write, avs_s1_writedata,
		  char_ram_q, font_rom_q)	
	  variable v: display_regs_type;
		variable clk_en: std_logic;
		variable font_address: std_logic_vector(14 downto 0);
    variable font_bit: std_logic;		
		
		procedure nextLine is
		begin
		  if r.cursor_y = ROW_NUM-1 then
			  v.scroll_y := r.scroll_y + 1;
				v.state := st_clear_row;
			else	
				v.cursor_x := (others => '0');
				v.cursor_y := r.cursor_y + 1;
			end if;			
		end procedure nextLine;	
	begin
		v := r;

		v.display_clk_cnt := r.display_clk_cnt + 1;
    clk_en := r.display_clk_cnt(r.display_clk_cnt'high);		
		
		char_ram_cmd.rd_address <= get_address(r.rd_ptr_x, r.rd_ptr_y, r.scroll_y);
		char_ram_cmd.wr_address <= get_address(r.cursor_x, r.cursor_y, r.scroll_y);
		char_ram_cmd.wr_data <= r.sym;
		char_ram_cmd.wr <= '0';
		font_address := (r.font_row & "00000000000");
		font_address := font_address + ("000" & r.font_col & "00000000") + ("0000000" & char_ram_q);
		font_rom_address <= font_address(14 downto 3);
		font_bit := font_rom_q(CONV_INTEGER(r.font_lsb));	
	
		if clk_en = '1' then
			if r.hcnt = tms.h_sync_end then
				v.hsync := '0';	
				
				if r.vcnt = tms.v_sync_end then
					v.vsync := '0';	
					v.cursor_cnt := r.cursor_cnt + 1;
				end if;	
				if r.vcnt = tms.v_blank_start then
					v.vblank := '1';
				elsif r.vcnt = tms.v_blank_end then
					v.vblank := '0';
				end if;	
				if r.vcnt = tms.v_size then	
					v.vcnt := (others => '0');
					v.vsync := '1';
				else
					v.vcnt := r.vcnt + 1;
				end if;		
			end if;	
			if r.hcnt = tms.h_blank_start then
				v.hblank := '1';
			elsif r.hcnt = tms.h_blank_end then
				v.hblank := '0';
			end if;	
	    if r.hcnt = tms.h_size then
				v.hcnt := (others => '0');
				v.hsync := '1';
			else	
	      v.hcnt := r.hcnt + 1;
	    end if;				
			
			v.font_lsb := font_address(2 downto 0);
			
			if r.hblank = '0' then
				if r.font_col = FONT_WIDTH-1 then
					v.font_col := (others => '0');
				else	
				  v.font_col := r.font_col + 1;
				end if;	
				if r.font_col = FONT_WIDTH-2 then
					if r.rd_ptr_x = COL_NUM - 1 then
				    if r.font_row = FONT_HEIGHT-1 then
					    v.font_row := (others => '0');
					    v.rd_ptr_y := r.rd_ptr_y + 1;
				    else	
				      v.font_row := r.font_row + 1;
				    end if;						
					end if;	
					v.rd_ptr_x := r.rd_ptr_x + 1;
				end if;	
			else	
				v.font_col := (others => '0'); 
				v.rd_ptr_x := (others => '0'); 
			end if;	
	
			if r.vblank = '1' then							
				v.font_row := (others => '0');
				v.rd_ptr_y := (others => '0');
			end if;	
			
			case r.state is
				when st_clear_screen =>
					char_ram_cmd.wr_data <= x"20";
					char_ram_cmd.wr <= '1';
					if r.cursor_x = COL_NUM-1 then
						v.cursor_x := (others => '0'); 
						if r.cursor_y = ROW_NUM-1 then
							v.cursor_y := (others => '0');
							v.state := st_idle;	
						else
						  v.cursor_y := r.cursor_y + 1;	
						end if;	 
					else
						v.cursor_x := r.cursor_x + 1;
					end if;	
				when st_clear_row =>
					char_ram_cmd.wr_data <= x"20";
					char_ram_cmd.wr <= '1';
					if r.cursor_x = COL_NUM-1 then
						v.cursor_x := (others => '0');
						v.state := st_idle;	
					else
						v.cursor_x := r.cursor_x + 1;					
					end if;					
				when st_idle =>
				  if r.sym_rdy = '1' then
						case r.sym is	 
							when x"09" =>
							  v.state := st_tab;
							when x"0D" =>
							  v.cursor_x := (others => '0');
							when x"0A" =>
								nextLine;
							when others =>
								char_ram_cmd.wr_data <= r.sym;
								char_ram_cmd.wr <= '1';						
								if r.cursor_x /= COL_NUM-1 then
								  v.cursor_x := r.cursor_x + 1;								
								else	
									nextLine;
								end if;	
						end case;
						v.sym_rdy := '0';
					end if;	
				when st_tab =>
					char_ram_cmd.wr_data <= x"20";
					char_ram_cmd.wr <= '1';
					if r.cursor_x /= COL_NUM-1 then
					  if r.cursor_x(2 downto 0) = "111" then
						  v.state := st_idle;
						else
							v.cursor_x := r.cursor_x + 1;
						end if;
					else
						nextLine;
					end if;	
					
			end case;	
		end if;  -- clk_en

		if r.rd_ptr_x = r.cursor_x and r.rd_ptr_y = r.cursor_y then
			if r.font_row = FONT_HEIGHT-1 or r.font_row = FONT_HEIGHT-2 then
        if BLINKED_CURSOR = 0 or r.cursor_cnt(r.cursor_cnt'high) = '1' then 
	        font_bit := '1';
        end if;	
			end if;
		end if;			
		
		if font_bit = '1' then
			v.rcolor := COLOR_FG.r;
			v.gcolor := COLOR_FG.g;
			v.bcolor := COLOR_FG.b;
		else
			v.rcolor := x"00";
			v.gcolor := x"00";
			v.bcolor := x"00";						
		end if;			
		
		-- Avalon Bus operations
		avs_s1_readdata <= (others => '0');
		if r.state = st_idle then
			avs_s1_readdata(0) <= '1';
		end if;	

	  if avs_s1_chipselect = '1' then
		  if avs_s1_write = '1' then
			  v.sym := avs_s1_writedata;
			  v.sym_rdy := '1'; -- not r.sym_rdy;
		  end if;	
	  end if;		
		
		next_r <= v;
	end process next_state_proc;	
	
	process(reset, clk)
	begin
		if reset = '1' then		
			r.state <= st_clear_screen;
			
		  r.display_clk_cnt <= (others => '0');
	    r.hcnt <= (others => '0');
	    r.vcnt <= (others => '0');
	    r.hblank <= '1';
	    r.hsync <= '1';
	    r.vblank <= '1';
	    r.vsync <= '1';			
			
			r.cursor_x <= (others => '0');
			r.cursor_y <= (others => '0');
			r.rd_ptr_x <= (others => '0');
			r.rd_ptr_y <= (others => '0');
			r.scroll_y <= (others => '0'); 
			r.sym_rdy <= '0';
			
	    r.rcolor <= (others => '0'); 
			r.gcolor <= (others => '0');
			r.bcolor <= (others => '0');
			
			r.cursor_cnt <= (others => '0');
			
			r.sym_rdy <= '0';
		elsif rising_edge(clk) then	
			r <= next_r;
		end if;		
	end process;	

	char_ram_proc: process(clk)
	begin
		if rising_edge(clk) then
			if char_ram_cmd.wr = '1' then
				char_ram(CONV_INTEGER(char_ram_cmd.wr_address)) <= char_ram_cmd.wr_data;
			end if;	
			char_ram_q <= char_ram(CONV_INTEGER(char_ram_cmd.rd_address));			
		end if;
	end process char_ram_proc;	

	font_rom_proc: process(clk)
	begin
		if rising_edge(clk) then
			if font_rom_address < FONT_SIZE then 
			  font_rom_q <= font_rom(CONV_INTEGER(font_rom_address));	
			else
				font_rom_q <= (others => 'X');
			end if;	
		end if;
	end process font_rom_proc;	
	
  process (reset, clk)
  begin
    if reset = '1' then
	    blank_del <= '0';
			blank_del2 <= '0';
			blank_del3 <= '0';
	  elsif rising_edge(clk) then
		  blank_del3 <= blank_del2; 
			blank_del2 <= blank_del;
			blank_del <= blank;
	  end if;	
  end process;	

	blank <= r.hblank or r.vblank;
	
  nRAMDAC_BLANK <= not blank_del2; 
  nRAMDAC_SYNC <= '0';
  RAMDAC_CLK <= not clk;	
	
	HSYNC <= r.hsync xor tms.h_sync_inv;
	VSYNC <= r.vsync xor tms.v_sync_inv; 

  RED <= r.rcolor; 
  GREEN <= r.gcolor;
  BLUE <= r.bcolor;	
	
--	dvi_out: process(reset, clk)
--	begin
--	  if falling_edge(clk) then
--		  DVI_DE <= not blank_del2;			
--			if display_clk_cnt(0) = '0' then
--			  DVI_D <= gcolor(3 downto 0) & bcolor;
--			else
--			  DVI_D <= rcolor & gcolor(7 downto 4);
--			end if;
--	  end if;
--	end process dvi_out;
	
--	DVI_CLK <= display_clk;
end behaviour;
